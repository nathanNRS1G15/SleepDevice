// projNiosII.v

// Generated using ACDS version 13.1 182 at 2018.07.13.16:39:00

`timescale 1 ps / 1 ps
module projNiosII (
		input  wire        clk_clk,                                 //                              clk.clk
		input  wire [7:0]  pio_switches_external_connection_export, // pio_switches_external_connection.export
		output wire [7:0]  pio_led_external_connection_export,      //      pio_led_external_connection.export
		output wire [11:0] dram_external_addr,                      //                    dram_external.addr
		output wire [1:0]  dram_external_ba,                        //                                 .ba
		output wire        dram_external_cas_n,                     //                                 .cas_n
		output wire        dram_external_cke,                       //                                 .cke
		output wire        dram_external_cs_n,                      //                                 .cs_n
		inout  wire [15:0] dram_external_dq,                        //                                 .dq
		output wire [1:0]  dram_external_dqm,                       //                                 .dqm
		output wire        dram_external_ras_n,                     //                                 .ras_n
		output wire        dram_external_we_n,                      //                                 .we_n
		output wire        altpll_0_c0_clk,                         //                      altpll_0_c0.clk
		input  wire        reset_reset_n,                           //                            reset.reset_n
		output wire [7:0]  pio_lcd_control_export,                  //                  pio_lcd_control.export
		output wire [7:0]  pio_lcd_data_export                      //                     pio_lcd_data.export
	);

	wire         altpll_0_c1_clk;                                              // altpll_0:c1 -> [irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:altpll_0_c1_clk, new_sdram_controller_0:clk, nios2_qsys_0:clk, onchip_memory2_0:clk, pio_LCD_control:clk, pio_LCD_data:clk, pio_LED:clk, pio_Switches:clk, rst_controller:clk, spi_master:clk, spi_slave:clk, timer_0:clk]
	wire         spi_master_external_sclk;                                     // spi_master:SCLK -> spi_slave:SCLK
	wire         spi_master_external_ss_n;                                     // spi_master:SS_n -> spi_slave:SS_n
	wire         spi_master_external_mosi;                                     // spi_master:MOSI -> spi_slave:MOSI
	wire         spi_slave_external_miso;                                      // spi_slave:MISO -> spi_master:MISO
	wire  [31:0] mm_interconnect_0_pio_lcd_control_s1_writedata;               // mm_interconnect_0:pio_LCD_control_s1_writedata -> pio_LCD_control:writedata
	wire   [1:0] mm_interconnect_0_pio_lcd_control_s1_address;                 // mm_interconnect_0:pio_LCD_control_s1_address -> pio_LCD_control:address
	wire         mm_interconnect_0_pio_lcd_control_s1_chipselect;              // mm_interconnect_0:pio_LCD_control_s1_chipselect -> pio_LCD_control:chipselect
	wire         mm_interconnect_0_pio_lcd_control_s1_write;                   // mm_interconnect_0:pio_LCD_control_s1_write -> pio_LCD_control:write_n
	wire  [31:0] mm_interconnect_0_pio_lcd_control_s1_readdata;                // pio_LCD_control:readdata -> mm_interconnect_0:pio_LCD_control_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_switches_s1_address;                    // mm_interconnect_0:pio_Switches_s1_address -> pio_Switches:address
	wire  [31:0] mm_interconnect_0_pio_switches_s1_readdata;                   // pio_Switches:readdata -> mm_interconnect_0:pio_Switches_s1_readdata
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_writedata;               // mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	wire   [1:0] mm_interconnect_0_altpll_0_pll_slave_address;                 // mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	wire         mm_interconnect_0_altpll_0_pll_slave_write;                   // mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	wire         mm_interconnect_0_altpll_0_pll_slave_read;                    // mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_readdata;                // altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	wire  [15:0] mm_interconnect_0_spi_master_spi_control_port_writedata;      // mm_interconnect_0:spi_master_spi_control_port_writedata -> spi_master:data_from_cpu
	wire   [2:0] mm_interconnect_0_spi_master_spi_control_port_address;        // mm_interconnect_0:spi_master_spi_control_port_address -> spi_master:mem_addr
	wire         mm_interconnect_0_spi_master_spi_control_port_chipselect;     // mm_interconnect_0:spi_master_spi_control_port_chipselect -> spi_master:spi_select
	wire         mm_interconnect_0_spi_master_spi_control_port_write;          // mm_interconnect_0:spi_master_spi_control_port_write -> spi_master:write_n
	wire         mm_interconnect_0_spi_master_spi_control_port_read;           // mm_interconnect_0:spi_master_spi_control_port_read -> spi_master:read_n
	wire  [15:0] mm_interconnect_0_spi_master_spi_control_port_readdata;       // spi_master:data_to_cpu -> mm_interconnect_0:spi_master_spi_control_port_readdata
	wire  [63:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;              // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire  [12:0] mm_interconnect_0_onchip_memory2_0_s1_address;                // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;             // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                  // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                  // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [63:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;               // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [7:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;             // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest; // nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata;   // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address;     // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write;       // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read;        // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata;    // nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess; // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable;  // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire         nios2_qsys_0_data_master_waitrequest;                         // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire  [31:0] nios2_qsys_0_data_master_writedata;                           // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [24:0] nios2_qsys_0_data_master_address;                             // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire         nios2_qsys_0_data_master_write;                               // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire         nios2_qsys_0_data_master_read;                                // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire  [31:0] nios2_qsys_0_data_master_readdata;                            // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_debugaccess;                         // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                          // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire  [15:0] mm_interconnect_0_spi_slave_spi_control_port_writedata;       // mm_interconnect_0:spi_slave_spi_control_port_writedata -> spi_slave:data_from_cpu
	wire   [2:0] mm_interconnect_0_spi_slave_spi_control_port_address;         // mm_interconnect_0:spi_slave_spi_control_port_address -> spi_slave:mem_addr
	wire         mm_interconnect_0_spi_slave_spi_control_port_chipselect;      // mm_interconnect_0:spi_slave_spi_control_port_chipselect -> spi_slave:spi_select
	wire         mm_interconnect_0_spi_slave_spi_control_port_write;           // mm_interconnect_0:spi_slave_spi_control_port_write -> spi_slave:write_n
	wire         mm_interconnect_0_spi_slave_spi_control_port_read;            // mm_interconnect_0:spi_slave_spi_control_port_read -> spi_slave:read_n
	wire  [15:0] mm_interconnect_0_spi_slave_spi_control_port_readdata;        // spi_slave:data_to_cpu -> mm_interconnect_0:spi_slave_spi_control_port_readdata
	wire         mm_interconnect_0_new_sdram_controller_0_s1_waitrequest;      // new_sdram_controller_0:za_waitrequest -> mm_interconnect_0:new_sdram_controller_0_s1_waitrequest
	wire  [15:0] mm_interconnect_0_new_sdram_controller_0_s1_writedata;        // mm_interconnect_0:new_sdram_controller_0_s1_writedata -> new_sdram_controller_0:az_data
	wire  [21:0] mm_interconnect_0_new_sdram_controller_0_s1_address;          // mm_interconnect_0:new_sdram_controller_0_s1_address -> new_sdram_controller_0:az_addr
	wire         mm_interconnect_0_new_sdram_controller_0_s1_chipselect;       // mm_interconnect_0:new_sdram_controller_0_s1_chipselect -> new_sdram_controller_0:az_cs
	wire         mm_interconnect_0_new_sdram_controller_0_s1_write;            // mm_interconnect_0:new_sdram_controller_0_s1_write -> new_sdram_controller_0:az_wr_n
	wire         mm_interconnect_0_new_sdram_controller_0_s1_read;             // mm_interconnect_0:new_sdram_controller_0_s1_read -> new_sdram_controller_0:az_rd_n
	wire  [15:0] mm_interconnect_0_new_sdram_controller_0_s1_readdata;         // new_sdram_controller_0:za_data -> mm_interconnect_0:new_sdram_controller_0_s1_readdata
	wire         mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid;    // new_sdram_controller_0:za_valid -> mm_interconnect_0:new_sdram_controller_0_s1_readdatavalid
	wire   [1:0] mm_interconnect_0_new_sdram_controller_0_s1_byteenable;       // mm_interconnect_0:new_sdram_controller_0_s1_byteenable -> new_sdram_controller_0:az_be_n
	wire  [31:0] mm_interconnect_0_pio_lcd_data_s1_writedata;                  // mm_interconnect_0:pio_LCD_data_s1_writedata -> pio_LCD_data:writedata
	wire   [1:0] mm_interconnect_0_pio_lcd_data_s1_address;                    // mm_interconnect_0:pio_LCD_data_s1_address -> pio_LCD_data:address
	wire         mm_interconnect_0_pio_lcd_data_s1_chipselect;                 // mm_interconnect_0:pio_LCD_data_s1_chipselect -> pio_LCD_data:chipselect
	wire         mm_interconnect_0_pio_lcd_data_s1_write;                      // mm_interconnect_0:pio_LCD_data_s1_write -> pio_LCD_data:write_n
	wire  [31:0] mm_interconnect_0_pio_lcd_data_s1_readdata;                   // pio_LCD_data:readdata -> mm_interconnect_0:pio_LCD_data_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_led_s1_writedata;                       // mm_interconnect_0:pio_LED_s1_writedata -> pio_LED:writedata
	wire   [1:0] mm_interconnect_0_pio_led_s1_address;                         // mm_interconnect_0:pio_LED_s1_address -> pio_LED:address
	wire         mm_interconnect_0_pio_led_s1_chipselect;                      // mm_interconnect_0:pio_LED_s1_chipselect -> pio_LED:chipselect
	wire         mm_interconnect_0_pio_led_s1_write;                           // mm_interconnect_0:pio_LED_s1_write -> pio_LED:write_n
	wire  [31:0] mm_interconnect_0_pio_led_s1_readdata;                        // pio_LED:readdata -> mm_interconnect_0:pio_LED_s1_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;  // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;     // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                       // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                         // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_chipselect;                      // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire         mm_interconnect_0_timer_0_s1_write;                           // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                        // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                  // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [24:0] nios2_qsys_0_instruction_master_address;                      // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                         // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                     // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         irq_mapper_receiver0_irq;                                     // timer_0:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                     // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                     // spi_master:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                     // spi_slave:irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                       // irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_qsys_0_reset_n_reset_bridge_in_reset_reset, new_sdram_controller_0:reset_n, nios2_qsys_0:reset_n, onchip_memory2_0:reset, pio_LCD_control:reset_n, pio_LCD_data:reset_n, pio_LED:reset_n, pio_Switches:reset_n, rst_translator:in_reset, spi_master:reset_n, spi_slave:reset_n, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [nios2_qsys_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_qsys_0_jtag_debug_module_reset_reset;                   // nios2_qsys_0:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                           // rst_controller_001:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]

	projNiosII_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (altpll_0_c1_clk),                                              //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                              //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                           //                          .reset_req
		.d_address                             (nios2_qsys_0_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                              // custom_instruction_master.readra
	);

	projNiosII_jtag_uart_0 jtag_uart_0 (
		.clk            (altpll_0_c1_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	projNiosII_timer_0 timer_0 (
		.clk        (altpll_0_c1_clk),                         //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                 //   irq.irq
	);

	projNiosII_pio_LED pio_led (
		.clk        (altpll_0_c1_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_pio_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_led_s1_readdata),   //                    .readdata
		.out_port   (pio_led_external_connection_export)       // external_connection.export
	);

	projNiosII_pio_Switches pio_switches (
		.clk      (altpll_0_c1_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_pio_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_switches_s1_readdata), //                    .readdata
		.in_port  (pio_switches_external_connection_export)     // external_connection.export
	);

	projNiosII_new_sdram_controller_0 new_sdram_controller_0 (
		.clk            (altpll_0_c1_clk),                                           //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                           // reset.reset_n
		.az_addr        (mm_interconnect_0_new_sdram_controller_0_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_new_sdram_controller_0_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_new_sdram_controller_0_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_new_sdram_controller_0_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_new_sdram_controller_0_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_new_sdram_controller_0_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_new_sdram_controller_0_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_new_sdram_controller_0_s1_waitrequest),   //      .waitrequest
		.zs_addr        (dram_external_addr),                                        //  wire.export
		.zs_ba          (dram_external_ba),                                          //      .export
		.zs_cas_n       (dram_external_cas_n),                                       //      .export
		.zs_cke         (dram_external_cke),                                         //      .export
		.zs_cs_n        (dram_external_cs_n),                                        //      .export
		.zs_dq          (dram_external_dq),                                          //      .export
		.zs_dqm         (dram_external_dqm),                                         //      .export
		.zs_ras_n       (dram_external_ras_n),                                       //      .export
		.zs_we_n        (dram_external_we_n)                                         //      .export
	);

	projNiosII_onchip_memory2_0 onchip_memory2_0 (
		.clk        (altpll_0_c1_clk),                                  //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //       .reset_req
	);

	projNiosII_altpll_0 altpll_0 (
		.clk       (clk_clk),                                        //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset),             // inclk_interface_reset.reset
		.read      (mm_interconnect_0_altpll_0_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_altpll_0_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_altpll_0_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_altpll_0_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_altpll_0_pll_slave_writedata), //                      .writedata
		.c0        (altpll_0_c0_clk),                                //                    c0.clk
		.c1        (altpll_0_c1_clk),                                //                    c1.clk
		.areset    (),                                               //        areset_conduit.export
		.locked    (),                                               //        locked_conduit.export
		.phasedone ()                                                //     phasedone_conduit.export
	);

	projNiosII_spi_master spi_master (
		.clk           (altpll_0_c1_clk),                                          //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                          //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_master_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_master_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_master_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_master_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_master_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_master_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver2_irq),                                 //              irq.irq
		.MISO          (spi_slave_external_miso),                                  //         external.export
		.MOSI          (spi_master_external_mosi),                                 //                 .export
		.SCLK          (spi_master_external_sclk),                                 //                 .export
		.SS_n          (spi_master_external_ss_n)                                  //                 .export
	);

	projNiosII_spi_slave spi_slave (
		.clk           (altpll_0_c1_clk),                                         //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                         //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_slave_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_slave_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_slave_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_slave_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_slave_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_slave_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver3_irq),                                //              irq.irq
		.MISO          (spi_slave_external_miso),                                 //         external.export
		.MOSI          (spi_master_external_mosi),                                //                 .export
		.SCLK          (spi_master_external_sclk),                                //                 .export
		.SS_n          (spi_master_external_ss_n)                                 //                 .export
	);

	projNiosII_pio_LED pio_lcd_data (
		.clk        (altpll_0_c1_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_pio_lcd_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_lcd_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_lcd_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_lcd_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_lcd_data_s1_readdata),   //                    .readdata
		.out_port   (pio_lcd_data_export)                           // external_connection.export
	);

	projNiosII_pio_LED pio_lcd_control (
		.clk        (altpll_0_c1_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_pio_lcd_control_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_lcd_control_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_lcd_control_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_lcd_control_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_lcd_control_s1_readdata),   //                    .readdata
		.out_port   (pio_lcd_control_export)                           // external_connection.export
	);

	projNiosII_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c1_clk                                            (altpll_0_c1_clk),                                              //                                          altpll_0_c1.clk
		.clk_0_clk_clk                                              (clk_clk),                                                      //                                            clk_0_clk.clk
		.altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                           // altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
		.nios2_qsys_0_reset_n_reset_bridge_in_reset_reset           (rst_controller_reset_out_reset),                               //           nios2_qsys_0_reset_n_reset_bridge_in_reset.reset
		.nios2_qsys_0_data_master_address                           (nios2_qsys_0_data_master_address),                             //                             nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest                       (nios2_qsys_0_data_master_waitrequest),                         //                                                     .waitrequest
		.nios2_qsys_0_data_master_byteenable                        (nios2_qsys_0_data_master_byteenable),                          //                                                     .byteenable
		.nios2_qsys_0_data_master_read                              (nios2_qsys_0_data_master_read),                                //                                                     .read
		.nios2_qsys_0_data_master_readdata                          (nios2_qsys_0_data_master_readdata),                            //                                                     .readdata
		.nios2_qsys_0_data_master_write                             (nios2_qsys_0_data_master_write),                               //                                                     .write
		.nios2_qsys_0_data_master_writedata                         (nios2_qsys_0_data_master_writedata),                           //                                                     .writedata
		.nios2_qsys_0_data_master_debugaccess                       (nios2_qsys_0_data_master_debugaccess),                         //                                                     .debugaccess
		.nios2_qsys_0_instruction_master_address                    (nios2_qsys_0_instruction_master_address),                      //                      nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest                (nios2_qsys_0_instruction_master_waitrequest),                  //                                                     .waitrequest
		.nios2_qsys_0_instruction_master_read                       (nios2_qsys_0_instruction_master_read),                         //                                                     .read
		.nios2_qsys_0_instruction_master_readdata                   (nios2_qsys_0_instruction_master_readdata),                     //                                                     .readdata
		.altpll_0_pll_slave_address                                 (mm_interconnect_0_altpll_0_pll_slave_address),                 //                                   altpll_0_pll_slave.address
		.altpll_0_pll_slave_write                                   (mm_interconnect_0_altpll_0_pll_slave_write),                   //                                                     .write
		.altpll_0_pll_slave_read                                    (mm_interconnect_0_altpll_0_pll_slave_read),                    //                                                     .read
		.altpll_0_pll_slave_readdata                                (mm_interconnect_0_altpll_0_pll_slave_readdata),                //                                                     .readdata
		.altpll_0_pll_slave_writedata                               (mm_interconnect_0_altpll_0_pll_slave_writedata),               //                                                     .writedata
		.jtag_uart_0_avalon_jtag_slave_address                      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),      //                        jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),        //                                                     .write
		.jtag_uart_0_avalon_jtag_slave_read                         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),         //                                                     .read
		.jtag_uart_0_avalon_jtag_slave_readdata                     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),     //                                                     .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),    //                                                     .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),  //                                                     .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),   //                                                     .chipselect
		.new_sdram_controller_0_s1_address                          (mm_interconnect_0_new_sdram_controller_0_s1_address),          //                            new_sdram_controller_0_s1.address
		.new_sdram_controller_0_s1_write                            (mm_interconnect_0_new_sdram_controller_0_s1_write),            //                                                     .write
		.new_sdram_controller_0_s1_read                             (mm_interconnect_0_new_sdram_controller_0_s1_read),             //                                                     .read
		.new_sdram_controller_0_s1_readdata                         (mm_interconnect_0_new_sdram_controller_0_s1_readdata),         //                                                     .readdata
		.new_sdram_controller_0_s1_writedata                        (mm_interconnect_0_new_sdram_controller_0_s1_writedata),        //                                                     .writedata
		.new_sdram_controller_0_s1_byteenable                       (mm_interconnect_0_new_sdram_controller_0_s1_byteenable),       //                                                     .byteenable
		.new_sdram_controller_0_s1_readdatavalid                    (mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid),    //                                                     .readdatavalid
		.new_sdram_controller_0_s1_waitrequest                      (mm_interconnect_0_new_sdram_controller_0_s1_waitrequest),      //                                                     .waitrequest
		.new_sdram_controller_0_s1_chipselect                       (mm_interconnect_0_new_sdram_controller_0_s1_chipselect),       //                                                     .chipselect
		.nios2_qsys_0_jtag_debug_module_address                     (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //                       nios2_qsys_0_jtag_debug_module.address
		.nios2_qsys_0_jtag_debug_module_write                       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                                                     .write
		.nios2_qsys_0_jtag_debug_module_read                        (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                                                     .read
		.nios2_qsys_0_jtag_debug_module_readdata                    (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                                                     .readdata
		.nios2_qsys_0_jtag_debug_module_writedata                   (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                                                     .writedata
		.nios2_qsys_0_jtag_debug_module_byteenable                  (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                                                     .byteenable
		.nios2_qsys_0_jtag_debug_module_waitrequest                 (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                                                     .waitrequest
		.nios2_qsys_0_jtag_debug_module_debugaccess                 (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                                                     .debugaccess
		.onchip_memory2_0_s1_address                                (mm_interconnect_0_onchip_memory2_0_s1_address),                //                                  onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                  (mm_interconnect_0_onchip_memory2_0_s1_write),                  //                                                     .write
		.onchip_memory2_0_s1_readdata                               (mm_interconnect_0_onchip_memory2_0_s1_readdata),               //                                                     .readdata
		.onchip_memory2_0_s1_writedata                              (mm_interconnect_0_onchip_memory2_0_s1_writedata),              //                                                     .writedata
		.onchip_memory2_0_s1_byteenable                             (mm_interconnect_0_onchip_memory2_0_s1_byteenable),             //                                                     .byteenable
		.onchip_memory2_0_s1_chipselect                             (mm_interconnect_0_onchip_memory2_0_s1_chipselect),             //                                                     .chipselect
		.onchip_memory2_0_s1_clken                                  (mm_interconnect_0_onchip_memory2_0_s1_clken),                  //                                                     .clken
		.pio_LCD_control_s1_address                                 (mm_interconnect_0_pio_lcd_control_s1_address),                 //                                   pio_LCD_control_s1.address
		.pio_LCD_control_s1_write                                   (mm_interconnect_0_pio_lcd_control_s1_write),                   //                                                     .write
		.pio_LCD_control_s1_readdata                                (mm_interconnect_0_pio_lcd_control_s1_readdata),                //                                                     .readdata
		.pio_LCD_control_s1_writedata                               (mm_interconnect_0_pio_lcd_control_s1_writedata),               //                                                     .writedata
		.pio_LCD_control_s1_chipselect                              (mm_interconnect_0_pio_lcd_control_s1_chipselect),              //                                                     .chipselect
		.pio_LCD_data_s1_address                                    (mm_interconnect_0_pio_lcd_data_s1_address),                    //                                      pio_LCD_data_s1.address
		.pio_LCD_data_s1_write                                      (mm_interconnect_0_pio_lcd_data_s1_write),                      //                                                     .write
		.pio_LCD_data_s1_readdata                                   (mm_interconnect_0_pio_lcd_data_s1_readdata),                   //                                                     .readdata
		.pio_LCD_data_s1_writedata                                  (mm_interconnect_0_pio_lcd_data_s1_writedata),                  //                                                     .writedata
		.pio_LCD_data_s1_chipselect                                 (mm_interconnect_0_pio_lcd_data_s1_chipselect),                 //                                                     .chipselect
		.pio_LED_s1_address                                         (mm_interconnect_0_pio_led_s1_address),                         //                                           pio_LED_s1.address
		.pio_LED_s1_write                                           (mm_interconnect_0_pio_led_s1_write),                           //                                                     .write
		.pio_LED_s1_readdata                                        (mm_interconnect_0_pio_led_s1_readdata),                        //                                                     .readdata
		.pio_LED_s1_writedata                                       (mm_interconnect_0_pio_led_s1_writedata),                       //                                                     .writedata
		.pio_LED_s1_chipselect                                      (mm_interconnect_0_pio_led_s1_chipselect),                      //                                                     .chipselect
		.pio_Switches_s1_address                                    (mm_interconnect_0_pio_switches_s1_address),                    //                                      pio_Switches_s1.address
		.pio_Switches_s1_readdata                                   (mm_interconnect_0_pio_switches_s1_readdata),                   //                                                     .readdata
		.spi_master_spi_control_port_address                        (mm_interconnect_0_spi_master_spi_control_port_address),        //                          spi_master_spi_control_port.address
		.spi_master_spi_control_port_write                          (mm_interconnect_0_spi_master_spi_control_port_write),          //                                                     .write
		.spi_master_spi_control_port_read                           (mm_interconnect_0_spi_master_spi_control_port_read),           //                                                     .read
		.spi_master_spi_control_port_readdata                       (mm_interconnect_0_spi_master_spi_control_port_readdata),       //                                                     .readdata
		.spi_master_spi_control_port_writedata                      (mm_interconnect_0_spi_master_spi_control_port_writedata),      //                                                     .writedata
		.spi_master_spi_control_port_chipselect                     (mm_interconnect_0_spi_master_spi_control_port_chipselect),     //                                                     .chipselect
		.spi_slave_spi_control_port_address                         (mm_interconnect_0_spi_slave_spi_control_port_address),         //                           spi_slave_spi_control_port.address
		.spi_slave_spi_control_port_write                           (mm_interconnect_0_spi_slave_spi_control_port_write),           //                                                     .write
		.spi_slave_spi_control_port_read                            (mm_interconnect_0_spi_slave_spi_control_port_read),            //                                                     .read
		.spi_slave_spi_control_port_readdata                        (mm_interconnect_0_spi_slave_spi_control_port_readdata),        //                                                     .readdata
		.spi_slave_spi_control_port_writedata                       (mm_interconnect_0_spi_slave_spi_control_port_writedata),       //                                                     .writedata
		.spi_slave_spi_control_port_chipselect                      (mm_interconnect_0_spi_slave_spi_control_port_chipselect),      //                                                     .chipselect
		.timer_0_s1_address                                         (mm_interconnect_0_timer_0_s1_address),                         //                                           timer_0_s1.address
		.timer_0_s1_write                                           (mm_interconnect_0_timer_0_s1_write),                           //                                                     .write
		.timer_0_s1_readdata                                        (mm_interconnect_0_timer_0_s1_readdata),                        //                                                     .readdata
		.timer_0_s1_writedata                                       (mm_interconnect_0_timer_0_s1_writedata),                       //                                                     .writedata
		.timer_0_s1_chipselect                                      (mm_interconnect_0_timer_0_s1_chipselect)                       //                                                     .chipselect
	);

	projNiosII_irq_mapper irq_mapper (
		.clk           (altpll_0_c1_clk),                //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                             // reset_in0.reset
		.reset_in1      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (altpll_0_c1_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),         //          .reset_req
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                             // reset_in0.reset
		.reset_in1      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                    //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

endmodule
